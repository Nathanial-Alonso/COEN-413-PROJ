`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GRDbaUVa+KMAvkCR4Jpxe50MvQ1gDfVSWHT/QbO9l1tJ/aoO5ojHUn7UVsENRI0y
oDFmt5wRuCRHvPqzPaAJhKtCBPR1Ea4LbO4r11fxHxBXN9NmHCYkVJg53nR2BeC3
UrEa8nUkA9DNkeXJRFMs5uYSyYJljaWmeH/hWcMnmcm4h7C8E6v/urt2OoZ2HrAn
VcXucmSfSBRmvO7uXu9gu0EKXg1QfhYvcMrJDKveUbn6E1CoNruJxHbiJxx937XW
fOWKc5+nj2wnCAUyyiUxEGGB/1I+lBqtl7dwgUacKE2QJdYeiyIuIt4pbMcqoJWf
0zBJpN7xFpzQxDFBnGK8Rn8jC6Vh4bUZwA20mokn1/6pGNajil8aHJUyEPGRrrvC
0ELlenUHDS82r3Erdo+wxnEAICtpdkQEkIhtvTutlLg5TpyXWhRRIt6V4k48Eof0
lFVdb94tPEJdnkFVhULPvMkVvjtmml2xpNJAnjvW7Pr3BD69uExbc3eHJGZ+EfUf
3PZjTvnoHQ7uMXK3kioWoMLL+FKqBfEloJ56uu82UbAFCa5xmIpp3OOADJsdnz/L
NsXBowHDUK/LXo1SesYpDm+DBdEbzt2tN4oq28+tikVqiupgVLld2i2G9QR+irMf
tgo5clRtOA8tdlyHcDd0QeZqBVsAFk0386SRbsx5riK3PsWFvw9fbQ21Ppr/6p33
0uVyYHFYFyL3rK3PBUHPj1aas+M6Byjp5Yvw0L+yv3RYAHTMUabU1zXEI+xHN2WH
8C3pFJ19nSlMs0NqaES38a6EKEOzx/0wb8+p4bCwVjspPrWCMdE1LO1aX8oCjGSa
Xsr5XtfHrTVsR+EFol3ha7HBR/KOwifcwg1NFC0X3+98OlI1GA3y23rYgs20n8sG
vZpD5gXzkrn7pqAKOJLocNTW4sAE/P8l5+puiEerW0IQGPvn10FclZN6JPO0KHnh
VB8jD1iZG3rAlnlRHDMb7f+KFjwuiPt1RvPlNchgw3bAXi0wC2j7FRLkbHLKVrJX
4Q9ciiyjIGc5hZm9HwXYLSOclGbGoc75t/4hrL20sLugWNcYJfqMWmk4uFlI61qF
xwOSXMbV4Xm5vHjohG6pGj1klGv6MPEBhxwoPm2JeTSm7OSwqG7uJi76IumTnV9s
2YGPUu8NMgY5LngM2xhtqgVzoo5SrUXCuA2Ua3T36QbSREuGEjxFfF7V8b5Rt5j1
dOYu9pHfxu2WXht1nMBsekjN0qzaU1eDezvL6cbgc+zR8hOqxX0BFl9NeLOoMnQL
8+hiWMiyXoJ3QYo+9HFBw96YNSF+CNB0M1L0a/gkF5gbhc9PBzfPGUyyVCSbihTQ
iZZt/lvN7aMWZrh/HGNV9p/lkrONRirazKz8Bgm+CTmliM9P9wuBPfMy+icGssG+
bhxOqaR+oAQksNz2XHzBm4+44zdVrv40TidRreb1yyfQ74U2g91QvYDmGkiqymag
IFFF39tkqoHr5tFlsnoTZQ==
`protect END_PROTECTED
