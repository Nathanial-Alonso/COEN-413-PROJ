`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KX/J238+XkoTzchnXrBjDLcxED/JvhB0v5DNYoXrl+eAyTsxEbb74MwhYKY9HDY4
8ei8/3L7ZMwSAkqUBfxsF2yVkWAI5ZooYgX/PJN52CWwxlE7rNKJf2daX3OWTvvu
IUbeX1lKyKHBRb4JqeQent7S76cssbPHJnsuEYTxXfvyoke9bpqhRUMifbs/fjY1
oAmL2mQaRwtR4EN/JNDmWVpCf2rmnM3GuuZdRuwAP/QSWf6tAq/SP182KJ9+c8W8
2Jdg2TRz0UeW22vVBIeh3cA0nlEGudeuplolfTxP429kDCCDq0C4qhx1nwns/+Bw
iaUkcoQRksafPAdfThTPGvZm34JaA0y2buT2flDUoPvuyAMNpBT7TSISuGof6f9d
HCQKvRpnPapsM8+ou1NAFxPpKCZ01NeEcmqsE9J9UVXbqjb1D5Ru1AkplIcXMvae
4753v4dhCNpOjE0M0X6SAIEuWMqj1En5FFgE7QU3OFNRnvMq8/HN1a4Wjeg4o/dA
6IT+1Uob8dCeh4yT1JsoUyYAB5bdAI0hYNSQLG9/R0xxTUafxc26AIjSY/blt3tu
I2bntGtfVpxEDSmV+OJWtHpTFZzqU+4OIomeoJQYw/HEgk90wDKVttBzTgcLRRhi
cnEw9CpwJQirE2lr1ILIeQ76dxD2JnSFHNbWgUoBk4KF3i1aFg2rytxY2tjTq1jT
GBRdyQjfbQafEsVGPb6d/4Fv38CpVGIwb8ft2rd9boJOMLXScrlkDoEZnQ98f1rY
w/QkEii65No31fiMXABSWtt3BzbWIqYRTbaDM8uCj3v6QtYMvmDIqgQtYIIugCK0
UOPWefjDbV32QY1bzz5HsMr+sG3rq44nigt7raVpAKXPRhvNTQj+P1UyK85GMp6G
tRz3zPD6J1rrMMfJM0x9XXZ/8xEijAcn8TUnN7dvdWSaMN5i9cK07bFJaX/vfoYV
vLk0VXXmj68bBol4uqhjrIRReVMgzCKfQBvCaoKK+s56KwCa0Jgvm/pY6RWCrQ1N
4ARhqiwzUzu7ceqEEncOv+tQlmNWs0Q1GRaxZ+wT88i4lWcRp2ptAiJClhi6fh0s
E7LmhVoDo9VrMgPl70f7WrcxdXpezUDQvhDjK8+UgNsgglvYMfH0eboFFE74o7kX
lseMuHG9fJFa6To1lbFjAniV009syzFWniaBrh4LfW2NTUA4oxXHLt5W8ji683Uw
k6ODOEULouWuQa8kJkKCsbDRf1wPsRQw8lkHGP+jLNzN9cSQDyryjQPuwvxXa5Y1
05f4BJ4bp2vFj/FgBZfwA6yf3sXXWuJa4mVfiDLwl/EYfrn20q/O4FvOXnEShvx+
qAV2U6QIHpc2UlAMLUNQS5vumx/vLv5ehrAlk/7+neIGGMOsX3BabivX+3wJHU05
J9A/Tn/900YzsPXQ75zzNGiNnItm9dEAa5WuPe4l8zC4+imaF9xjpi6VXYKQWWoT
uMFfcHWs0RF1lafXyCKmfMlDVO3g0rc2IXWAU5WHV9tVZ/MYDv1c+ZqJwBXf3VBL
pw4rFQUX3zoYCAg3jhPjBDc6FpFokapDE/nfCOEDF2u0KDcDV8ft7JAAESzJ3Jd3
lM92GsmgDUlYqjHuaUj8EwBS7MZ8s9/LxVXckiIUMhC87YcTFX7PLlb2RbaJX1JQ
B5foiySLhwYrnka9YrYmGWkUmU6cuK+qINbyrH0eaQZxEf5J25IKO/yXwSiMKIZ1
uu4jwxlQtSvsXqI0AU9mkup5V2KnL/43CyibEyTg6zXkOgp0Ct6aGZWsvMjYRl4e
Ai9fj4faP65irfhFPl5NF1sTrc0O8G5dcaL31lSdtO45Gy1Y3SygtxUR7kMyrFME
`protect END_PROTECTED
