`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9CXfvCZOAbE10T3RILniMXDSkKxuualJWW3gCWxHTAl00xmZcmXiz88SUBjzIqpH
R6pR8ndQNqhGlqfiQq56m80GTcbHRRbkykfzYZqJlYf64EaXUJRGyBj5EB6blpgK
8A6V/r3D14IlRqALhxLzMvEeYwGN5a31728PzzxQXTbv706h4zaO8KuhgSxSrshC
bNfQqfOzDpGtMHNSzIgepGQm7i4jEWpU8HCC6BN+81sTQwXqgfM9NoItMtzBDBV6
VMyF+3LeyL8EPxkArc48qoc/Fpfm7O68eB57IdFV7JTyKrFB/yEtn6Gt3VbmsSkb
knOPeVgzJTQ4GPAkc01k5GjzIyh/G9EdwouxZiNBhmyzjYdE13ZemTvAzylxHR0W
zUDITaJqW0giuNiD71EFfc0k+6Cc7FuedydtB+9DJhLN4Er4+MGQ/5tt6Pb7zUUE
HU+vvCqNJXi4YUq5lNxSs1Uc9emRd0pYBWz/+C7Eh5ZTdvxGKiNGYqd5x9/6xu7Q
fm2eWXP03quQQcO27qZjWdpBsKcZRNKSL4u3tOTDoeRoCpt5pxd/X1Ho30wmni4R
140AmVD76LavpBlVIZVMJT7dBlvJk6an+ToVceC9Qzpo58cI5ZmQcoQXV6zhoAcF
YMAa6uI6PjU63AQpHnHjmlbN6IineGt0V9tsz6oWRZL2iHH5969MKivx4rdHlCRd
Jg9HSi4TazmeN5Hx0R/mQ4YoE/gDAsvU7sLMejzAKFr5kVwkw8MyJrRScMixSSdO
DB12pjVP33tDM1aGP0+/TnLcKHMkUmjrvA3YMJJWqEnxT4gb+ZUgaWuTFicBDwrV
QXDvkBpRZ1Bdd8+bMbJx5skZmRUlR5tETWM2oCxepsak5TRU72UkOpl7hrb4680S
o3vTxTJeuhqcb8ny9KXTWKpya294CXnebzdWsKEDOp5uBY4kQWsjnlsPFmH1I1cn
erQnEAWxVlVHLSl7MH6Sr9orRey46WROrtC4ZYb7jmvh+M5G5cZoj0OU7hc8licp
y9YvMbR0m4Tae2B4nBcmSSSlyGpHxfTKI/KbUjZ+Btf/MICPVMXNZz+el9FK6x1f
npYMvEan82XgEF/8QPW/u8lxs5duWeXLpLezHJUZ9n+SuovGJa0Snnxbxa/WvukE
n/+rb4QFqbyQQ/su3PBf35TmFUPsBYHdrrxZSPHuUZ5aVczvFRW/hwQi+rhVUBzc
Ow3CWPMW9iFx1caGxFLuXA1DnruuvM/5/MTisvSTS+ujBUsp4Z8ApMQo+yHphlaO
BxEYS4qPawzShX3m3N7dlhDunSiw+PL1V5h50LpMXfIhlgIvLT3SO/akVaGp525L
jwycJo8+OiF10PEzmJ7hGlmoQWtPGYQWzvjZECZVWyf4aj05KeGJCwG4MSLE5WX5
aRvvRyAovOGvA7Klfk8Ahs53iUFDYORYD1hBe0bSaccv/UF32GLO45U0rILAhFCe
gYEptraUInfn6uKVqeVbrg==
`protect END_PROTECTED
