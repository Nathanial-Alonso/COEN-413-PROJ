`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZV5JYhSw/5wzvqBN+kXQz298OVn7iZMFDDJUk/GAJUW4KjWQE1salTLbse4DCQy
t6hZeGvqX9ERS+vKxMcxg6dN+t/o2OCTwu/B6PMNUcYtsqVYHDPFmWa7C7Q9DXNW
E1GquobrO2Kr0aoN76Qdakmj4ZzT3+IQs0BJuzW561vmTPKom7Vc5a9F5cgRCt4O
Zv1bwmtI9gbfO3tr1xwmqhmK8meSYSHa8gIxrXjhRdPeFyulMKXeIDt+deu/7HEF
+lGXt0KNg6OPnKxAeqdkYMOP6K7kirbRNU/O+HUjDDAAPNWqCPi0KCN9n9F6degm
AiPqvKeKrfvpCvnDk4KGmGlHlx8ngcp6FtixN6dj8GFsp/52mqYU7cJqsRy/Pja6
ZtjlMR5XNcZVY3TIhgmewlqp4nyQs0QGJI7/BcBaz19fRO/jhDL0C2IyupaqILHb
mTn66wTbaY86bmEnsBGOh/IVcXFyOLQBmN/xLRcsRfz/9rsCoRVvHZq3lDbMtbqx
lc4Snj3D9jxU+UafuV+B/lge1exdlOGTkBoI6K1Xl7Y1UzQFhNgI2Nc6ZhE9H5mb
/ufMAVDuQ6+E8DhdvwtcaplJFzDLbH6h6MvslBNkGcRzTja89vOerD0NPfW+58O8
vKFKDRYhmvM5hITiYOf2sTyyxxZAZ7AonIX9jT86GmuT0Humt/OHtVVw49fedfQx
iloQUDVfijjE9LGFLzvNd8IkCcPQjkA6dRGZYUIgkqyHuBvN2cUiOpcJ9tOxKC/K
u3VomuTAd4pm1ixOQl9ram3HAgU+cImcTsCFUC1yditraHZ6k6wLdV6q/HjnFfcM
OZPLFn1xz8lwFKsdG+6Sc8bdC/Hn6s1HVTbjHwePOVUFguAaB0CqDl1yI0qERshh
HpH9BpFiIVo4T2/oYMlsPskZ9w43R83RsJrhqAP0TYQXB1dvDKR3Borne4RcyEHW
dEqy/0A1j0wlzX6Htxv94tBqBlxi/Sfvmx1tBg7hBFGy2bJ4rMuQPrprqvxheBIW
o+dWgE6MCUnMU/PdJuY8BEwY0/2Loj2+ACnrmjnlyoF/9EXYKm7DXCXpN4EX1+rH
FVHUwr/V76PnYQpR6LZVrw==
`protect END_PROTECTED
