`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FovBAlbC60l6fI0TL86JcKbVAQvmpyHAxN54ywDiuDplxRWCF1k/2IzV/LyN3az0
kbeTegftNBupaSOLgq297Du0jnHwfEb2cvS1BHM8xmtjIjauOXK/+C9V8bB7cTKI
1mb+s6Tp3x8KniQd2mFvG+FlUUJScN17Rs0D5R01zatu3Kg2XdrcXxyGTXC0i58n
1FBrAYTQSOQKfygxKKWUzyUHWAqL6J7n4J8jG0JZPE6Jam18xba5RNJfNsMdI5ON
wRtxeECjSQut2kEpvl/zoKfh1wXWYp8SexP/AOEOmFT7X1sN4YhhY8jX70ykaUE8
ekwwaVUMZ51l41uyk9hji+SdMcjKGWfeF5uA8bHd/3LlXxrm3+1i1gGfBehS501r
+0GYZme86SG9/eujXXhSRbqSHipYmhoa5DgR4GqLPOxkzCdxdFUkDgwyG2iOaWaB
rZwv2YZt1aHsUGSGrh1Xjn7KpdEP6Y4aVsB4ButpyqaOlCA7vV43Yg+mudER9Z8t
kqqj+rda2HkYSzk/oWi/f6bR5yN3BKHQWCAp1KNW4nT1n/z16qP+N/fVv7z/Su1U
`protect END_PROTECTED
