`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mVE8P4rayCyud6Z1pAH79E8NOYi1Y7kBrP717LNpPyUxhNLQFI1mWy5TXF9uqnYi
CR+QbfDghr2SZWKZyxP41OOMJjk2GePCKEi95um5LOR4cl7inm7MuMtzE48tkXIP
w5JYrxxMvhAQHG9axU0ACBGp2t0fG41pW6OkNyXaJNnYweoISvVT30T9TkcI8Grp
dU1i5HSMNpTuUGQ80Zeh+Hb4zJTnneacnqhokk17r9pILmcheb2mQxM6CME2rO6M
7eA8OzdzgAHqmPehke+E+/kVGCWSMDPsyC5icvxrd0vKvnjUQfybjo4HYwekOQNx
CrkIJhuO4Ukm0tg4neNQ6BpGAbULHcHv/vNzveossVIw1IAz/S+M0+/8amL5Lg/9
eLErrM/Buk1727irbujX2U7e5MmUo3aq/9DmMesjAsBoXgyToP80I+6gXkLObYdB
SEPwzWCmMUNEXzeR9/z0zzjbs6f3cSqB/tjbX6/cYXzrgmhJNNaK+Z0fudV2pw/j
1z01XCQWyDk4bgUJO6LNIIe0A+2o2Qzruc5abT9VYPSbvjLzfvjZZTp3ur0IJ6+1
kRYMgdSIwHdQDxhIgwVEKQ==
`protect END_PROTECTED
