`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JrFX7KPvCHGk7trz6yrj+dS625Q3lnbsx8KMJbAS7SoNNcWhGlSLckr8fosOg7Zr
jy1EaJIKZIdenppMqbaSaTET+9fcbrfTBmUGCAEwu3SL142TvNYG7TquJ9QiRMUD
kVD2UIAB0yLZ5Cblfg6ywe1i7j0RFufnK3IjBRhEHXDczUtkrRStIYU8n0cm6wy+
H/NqIKcDHEsmOGJBDxFc4QCPINqBmzPyEkMFrfKfb/Jr3xTkABDKjaMygAv9nEz5
7rWpVeXQikhOFkgynjJMQjhDuwcjDCgV4kTwgiME95HELUPY5BrsUxuNYGfAWWQz
iPL7UrFSjsnXo2ogOEubkcN1SDEemmmZXt+clwyOwH1kNGyRSr9XS4mH/AGWLBti
a987nBb1/Jqs/bThT1hIDJptIJPAxafvhLn06jzATbrP7S2YhcbzXO/OCvPumlq2
+lqBuAgD6hW1KUrqe/CU4pkLJ17OIvXVEM8O2cF1Y3wlQz/fZFTkiEHD1S4z55cV
C90OVWg7YwHqzpuaWjLCHG6K/xCyNJ7c7+8hQzZHHWUPm3n3Z/9SLkWOW0vxa+eY
3wwdJXKkxkAYV9GKn/7XKGjNU9c+wfqK4f5yyKBkrTaNoGVB09KOtxn91eQFtKaz
z8vMbwNAcVgtWNnkk2B+9dyn3M7KbHwkIs/hOeu68r36qKZET7HUGS0zdPBtI7e1
jt09uW48zrNTNW9M7Z2lQ0jlGOQffpv6XWIXkPt0A7bGh8djuSWWwfeUVSuKPE/7
9XueXGo3CfgyEpP0dWWWIndcHR5apd8tyx4/gTqIjfa3AOUgh5SpbaeyV9Aw+oF4
v9BkD7UM1IpK93kfOjJcGQx878WizGX0GWOjpaRExWmvoDfMpaUFuT00M0suFDvS
6pyrnP6crOwAIYJ+hic+RA==
`protect END_PROTECTED
