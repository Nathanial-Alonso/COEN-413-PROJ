`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4orJxqR4dYzxpBxfC01tirMm1XmWGqFhMS2d2GLYxyjO6okw/07vLdOywOEQW9B8
+aOWfulxV7vTU7IAFB8X+en3GnDPO42fqI6yf8jP9Ul4qHsXbSQHOgWBSMw2sIEB
tOBEXupfwdtweurQkwM+oy8oix94CzUFg/Gh3k0P9ScuNd/+yWuMYbdJgp+DzSsL
CR+WA7CXUcqYYYq0qbS3qxikk0gGcznG1TUuo29rnlNuyTyEQ6d8NlLjvyuzxVrz
zN2xNAa7oyFHJubs1/mwNbRugYf3s4SKnZOLWGzLeVtOTQIkCqbWc2QtOG5YOq81
qaHblr1HyS08FKJdxue+25LLy3r8IHfob/WiEYF1FQx4cQ9gVxte5fzll2T0TieD
7A6vOneEWUhpuPGnH0ctneC8R4qRWwMBQiyUvUgXxGG22LzTK+BHwDZ3EbxTNoVh
Sw76ov41FqEJC94kZ0PW1umFbGW7KzCZiSALmBXjKpADOa8c3sBaxD+oF/kY9l/3
fCmgxmB9e5AdM5H64uVRFYu446KiI/U7/NqrwuaM7uGkZ3doML3emfmPh2wFuX71
VL0NkHGI3f0xudRmkU4XzUwegwvxdcoHM5znebRRRDI=
`protect END_PROTECTED
