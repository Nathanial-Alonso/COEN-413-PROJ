library verilog;
use verilog.vl_types.all;
entity TestTop is
end TestTop;
