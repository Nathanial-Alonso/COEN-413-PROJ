library verilog;
use verilog.vl_types.all;
entity calcInterface is
    port(
        clk             : in     vl_logic
    );
end calcInterface;
