program test(dut_if IF);
 import classes::*;
 Generator generator;
 Agent agent;
 Scoreboard scoreboard;
 Checker checker;
 Driver driver;
 Monitor monitor;


 inital begin
     
 

 end

endprogram

